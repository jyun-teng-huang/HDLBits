module top_module (
    input a,
    input b,
    output q );//

    assign q = b&a; // Fix me

endmodule
